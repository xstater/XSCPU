`ifndef _RAM_VH_
`define _RAM_VH_

`include "src/defs.vh"

`define RAM_SIZE 128
`define RAM_ADDR_WIDTH 8:0
`define RAM_DATA_WIDTH 31:0

`define RAM_WRITE 1'b1
`define RAM_READ  1'b0

`endif