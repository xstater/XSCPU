`ifndef _PC_H_
`define _PC_H_

`include "src/defs.vh"

`define PC_ADDR_WIDTH 32
`define PC_ADDR_WIDTH_VECTOR (`PC_ADDR_WIDTH-1):0


`endif 