`ifndef _DEFS_H_
`define _DEFS_H_

`default_nettype none

`define HIGH 1'b1
`define LOW  1'b0
`define ENABLE  1'b1
`define DISABLE 1'b0


`endif //_DEFS_H_